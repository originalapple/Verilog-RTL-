always @*
begin
    out1 = a? b+c:d+e;
    out2 = f? g+h:p+m;

end
